module gf180mcu_name_plate;
endmodule
